//Define package and include all files
package apb_pkg;
`include "uvm_macros.svh"
 import uvm_pkg::*;
	`include "apb_master_config.sv"
  `include "apb_slave_config.sv"
  `include "apb_base_seq_item.sv"
	`include "apb_master_seq.sv"
	`include "apb_slave_seq.sv"
	`include "apb_master_sequencer.sv"
	`include "apb_slave_sequencer.sv"
	`include "apb_master_driver.sv"
	`include "apb_master_monitor.sv"
	`include "apb_master_agent.sv"
	`include "apb_slave_driver.sv"
	`include "apb_slave_monitor.sv"
	`include "apb_slave_agent.sv"
  `include "apb_virtual_sequencer.sv"
endpackage
